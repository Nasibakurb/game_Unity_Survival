    ����          Assembly-CSharp   SaveGame+Position   xyz      ǽEǽEǽE